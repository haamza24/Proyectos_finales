library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity programa_helloworld_int_FLIP is
	port( address : in std_logic_vector(7 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(15 downto 0));
	end;

architecture v1 of programa_helloworld_int_FLIP is

	constant ROM_WIDTH: INTEGER:= 16;
	constant ROM_LENGTH: INTEGER:= 256;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"1111000000000000",
	"1101100011001100",
	"1000101001000111",
	"0100000101000000",
	"1101100011011001",
	"0100000001000000",
	"0011001000101010",
	"1101010100100110",
	"1101100000101111",
	"1101100011001100",
	"1000101001000001",
	"0100000101000000",
	"1101100011011001",
	"1101100011001100",
	"1000101001000010",
	"0100000101000000",
	"1101100011011001",
	"1101100010010100",
	"1101100010010100",
	"1101100001100011",
	"1101100011001100",
	"1000101001000011",
	"0100000101000000",
	"1101100011011001",
	"1101100011001100",
	"1000101001000100",
	"0100000101000000",
	"1101100011011001",
	"1101100011001100",
	"1000101001000100",
	"0100000101000000",
	"1101100011011001",
	"1101100010010100",
	"1101100010011011",
	"1000000101010000",
	"1101100011011001",
	"1101100010010100",
	"1101000000000001",
	"0011000001110010",
	"1101010100100110",
	"1000000101100001",
	"1000100101000001",
	"1101100011011001",
	"1000000101100010",
	"1000100101000010",
	"1101100011011001",
	"1101100000010010",
	"0000000001001001",
	"0100000100000000",
	"1101100011011001",
	"0000000001101110",
	"0100000100000000",
	"1101100011011001",
	"0000000001110100",
	"0100000100000000",
	"1101100011011001",
	"0000000001110010",
	"0100000100000000",
	"1101100011011001",
	"0000000001101111",
	"0100000100000000",
	"1101100011011001",
	"0000000001100100",
	"0100000100000000",
	"1101100011011001",
	"0000000001110101",
	"0100000100000000",
	"1101100011011001",
	"0000000001100011",
	"0100000100000000",
	"1101100011011001",
	"0000000001100101",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"0000000001100011",
	"0100000100000000",
	"1101100011011001",
	"0000000001101100",
	"0100000100000000",
	"1101100011011001",
	"0000000001100001",
	"0100000100000000",
	"1101100011011001",
	"0000000001110110",
	"0100000100000000",
	"1101100011011001",
	"0000000001100101",
	"0100000100000000",
	"1101100011011001",
	"0000000000111010",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"1001000000000000",
	"0000000001001001",
	"0100000100000000",
	"1101100011011001",
	"0000000001101110",
	"0100000100000000",
	"1101100011011001",
	"0000000001110100",
	"0100000100000000",
	"1101100011011001",
	"0000000001110010",
	"0100000100000000",
	"1101100011011001",
	"0000000001101111",
	"0100000100000000",
	"1101100011011001",
	"0000000001100100",
	"0100000100000000",
	"1101100011011001",
	"0000000001110101",
	"0100000100000000",
	"1101100011011001",
	"0000000001100011",
	"0100000100000000",
	"1101100011011001",
	"0000000001100101",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"0000000001100100",
	"0100000100000000",
	"1101100011011001",
	"0000000001100001",
	"0100000100000000",
	"1101100011011001",
	"0000000001110100",
	"0100000100000000",
	"1101100011011001",
	"0000000001101111",
	"0100000100000000",
	"1101100011011001",
	"0000000000111010",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"1001000000000000",
	"0000000000001010",
	"0100000100000000",
	"1101100011011001",
	"0000000000001101",
	"0100000100000000",
	"1101100011011001",
	"1001000000000000",
	"0000000001010100",
	"0100000100000000",
	"1101100011011001",
	"0000000001110101",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"0000000001100100",
	"0100000100000000",
	"1101100011011001",
	"0000000001100001",
	"0100000100000000",
	"1101100011011001",
	"0000000001110100",
	"0100000100000000",
	"1101100011011001",
	"0000000001101111",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"0000000001100101",
	"0100000100000000",
	"1101100011011001",
	"0000000001110011",
	"0100000100000000",
	"1101100011011001",
	"0000000000111010",
	"0100000100000000",
	"1101100011011001",
	"0000000000100000",
	"0100000100000000",
	"1101100011011001",
	"1001000000000000",
	"1100000111100000",
	"0010000100000000",
	"1101010011000110",
	"1101100011011001",
	"0010011100000001",
	"1101000011000000",
	"1111000000000001",
	"0000011000001001",
	"0011011000000001",
	"1101010111001000",
	"0000011000001001",
	"1101000011001000",
	"1000001011111111",
	"0000101010000000",
	"1101010111001100",
	"1101100011101101",
	"0000001100001001",
	"1101100011100110",
	"1010001000001110",
	"1000000011111111",
	"0000100010000000",
	"0101001000000000",
	"0011001100000001",
	"1101010111010001",
	"1001000000000000",
	"0000000000000000",
	"1000100011111111",
	"1101100011100110",
	"0000001100001000",
	"1000100111111111",
	"1101100011100110",
	"1010000100001110",
	"0011001100000001",
	"1101010111011101",
	"0000000011111111",
	"1000100011111111",
	"1101100011100110",
	"1001000000000000",
	"0000010000000011",
	"0000010100100010",
	"0011010100000001",
	"1101010111101000",
	"0011010000000001",
	"1101010111100111",
	"1001000000000000",
	"0000010000000011",
	"0000010100010000",
	"0011010100000001",
	"1101010111101111",
	"0011010000000001",
	"1101010111101110",
	"1001000000000000",
	"1111000000000000",
	"1101100011001100",
	"1111101000000000",
	"0100000101000000",
	"1101100011011001",
	"0010011000110000",
	"0100000111000000",
	"1101100011011001",
	"1011000000000001",
	"0000000000000000",
	"0000000000000000",
	"1101000011110100");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
